----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:30:06 04/20/2017 
-- Design Name: 
-- Module Name:    hx711 - a_hx711 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity hx711 is
	port( clk : in std_logic;
			DOUT: in std_logic;			--data from the hx711 module(24 bits, one by one starting with the MSB)
			SCK: out std_logic;		--clock generated by us with a frequency of 500KHz (T = 2 us)
			an: out std_logic_vector(3 downto 0);
			cat: out std_logic_vector(6 downto 0);
			dp: out std_logic;
			led: out std_logic_vector(7 downto 0));
end hx711;


architecture a_hx711 of hx711 is

component seven_seg is
	port(seg3, seg2, seg1, seg0: in std_logic_vector(3 downto 0);
			clk: in std_logic;
			an: out std_logic_vector(3 downto 0);
			cat: out std_logic_vector(6 downto 0));
end component;

signal seven_seg3, seven_seg2, seven_seg1, seven_seg0: std_logic_vector(3 downto 0); --the 4 seven segment displays

type states is (INIT, START, WAIT_BEFORE_READ, READ_DATA);
signal state: states;

signal count_wait: std_logic_vector(2 downto 0) := (others => '0');
signal count_read: std_logic_vector(11 downto 0) := (others => '0'); --count to 2500 (25 * 100 ns == 25 * ( 50 high + 50 low))

signal data, final_data : std_logic_vector(23 downto 0);
signal shift: std_logic := '0';

signal en_cnt_50, rst_cnt_50: std_logic := '0';
signal clock_500KHz: std_logic :=  '0';
signal count_50 : std_logic_vector(5 downto 0) := (others => '0');

signal falling_edge_500KHz: std_logic_vector(1 downto 0) := (others => '0');
begin

	
	DISPLAY: seven_seg port map (seven_seg3, seven_seg2, seven_seg1, seven_seg0, clk, an, cat);
	
	process(clk, final_data)
	begin
		if rising_edge(clk) then
			led <= final_data(23 downto 16);--most significant 8 bits
			seven_seg3 <= final_data(15 downto 12);
			seven_seg2 <= final_data(11 downto 8);
			seven_seg1 <= final_data(7 downto 4);
			seven_seg0 <= final_data(3 downto 0);
		end if;
	end process;
	
	process(clk, state, DOUT)
	begin
		if rising_edge(clk) then
			rst_cnt_50 <= '0';
			en_cnt_50 <= '0';
			
			case state is
				when INIT => if DOUT = '0' then
									state <= START;
								else
									state <= INIT;
								end if;
								
				when START => if DOUT = '0' then 
									state <= WAIT_BEFORE_READ;
								  else
									state <= INIT;	
								  end if;
								  
				when WAIT_BEFORE_READ => if DOUT = '1' then -- error => DOUT should be LOW 
													state <= INIT;
												 elsif count_wait = "101" then 
													state <= READ_DATA;
													count_wait <= (others => '0');
												 else
													state <= WAIT_BEFORE_READ;
													count_wait <= count_wait + 1;
												 end if;
												
	         when READ_DATA => if count_read = "100111000100" then --if count_read = 2500
											state <= INIT;
											final_data <= data ;--- x"FEA700";--pune intr o memorie o referinta < decat ceva
											count_read <= (others => '0');
											rst_cnt_50 <= '1';
										else
											state <= READ_DATA;
											count_read <= count_read + 1;
											en_cnt_50 <= '1';
										end if;
			end case;
		end if;
	end process;
	
	
	process(state, clock_500KHz)
	begin
		case state is
			when INIT => shift <= '0';
							 SCK <= '0';
			when START => shift <= '0';
							  SCK <= '0';
			when WAIT_BEFORE_READ => shift <= '0';
											 SCK <= '0';
			when READ_DATA => shift <= '1';
									SCK <= clock_500KHz;
		end case;
	end process;


	
	process(clk, en_cnt_50, rst_cnt_50, count_50, clock_500KHz)
	begin
	if rst_cnt_50 = '1' then
		count_50 <= (others => '0');-- counter will have the value 1
		clock_500KHz <= '0';
		falling_edge_500KHz <= (others => '0');
		
	elsif rising_edge(clk) then
			if en_cnt_50 = '1' then
				if count_50 = "110010" then -- if counter = 50
					count_50 <= "000001";-- counter will have the value 1
					
					if clock_500KHz = '1' then
						falling_edge_500KHz <= '1' & falling_edge_500KHz(1);
					else
						falling_edge_500KHz <= '0' & falling_edge_500KHz(1);
					end if;
					
					clock_500KHz <= not clock_500KHz;
					
				else
					falling_edge_500KHz <= '0' & falling_edge_500KHz(1);
					count_50 <= count_50 + 1;
				end if;
			end if;
	end if;
	end process;
	
	
	process(clk, shift, falling_edge_500KHz, DOUT)
	begin
		if rising_edge(clk) then
			if shift = '1' and falling_edge_500KHz = "10" then
				data <= data(22 downto 0) & DOUT;
			end if;
		end if;
	end process;
	
	dp <= '1';
end a_hx711;